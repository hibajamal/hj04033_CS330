module top(
  input [31:0] instruction,
  output reg [63:0] ReadData1,
  output reg [63:0] ReadData2
);